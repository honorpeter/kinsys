`ifndef _NINJIN_SVH_
`define _NINJIN_SVH_

`timescale 1 ns / 1 ps

package gobou;
  `include "gobou.svh"
endpackage

package renkon;
  `include "renkon.svh"
endpackage

`endif
