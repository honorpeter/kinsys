`ifndef _COMMON_SVH_
`define _COMMON_SVH_

`default_nettype wire
`timescale 1 ns / 1 ps
`define DIST

parameter STEP    = 10;
parameter DWIDTH  = 16;
parameter LWIDTH  = 10;
parameter IMGSIZE = 12;

parameter D_BIAS     = 2;
parameter D_RELU     = 2;

`endif
