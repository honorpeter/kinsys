module accum
endmodule
