`include "renkon.svh"

module renkon_ctrl_linebuf
 #(
  )
  ( input clk
  , input xrst
  );

endmodule
