`ifndef _NINJIN_SVH_
`define _NINJIN_SVH_

`include "common.svh"
`include "gobou.svh"
`include "renkon.svh"

parameter PORT = 32;

`endif
