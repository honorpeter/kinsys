`include "renkon.svh"

module renkon_ctrl_linebuf_pad
 #(
  )
  ( input clk
  , input xrst
  );

endmodule
