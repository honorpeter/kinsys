`ifndef _NINJIN_SVH_
`define _NINJIN_SVH_

`include "common.svh"

parameter PORT  = 32;
parameter LSB   = 2;

parameter ID_WIDTH      = 12;
parameter AWUSER_WIDTH  = 0;
parameter ARUSER_WIDTH  = 0;
parameter WUSER_WIDTH   = 0;
parameter RUSER_WIDTH   = 0;
parameter BUSER_WIDTH   = 0;

`endif
