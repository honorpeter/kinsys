parameter DWIDTH = 16;
parameter LWIDTH = 10;
parameter CORE   = 8;
parameter STEP   = 10;
