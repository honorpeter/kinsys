`include "renkon.svh"

module core
  (
  );

  conv conv(.*);

  bias bias(.*);

  relu relu(.*);

  pool pool(.*);

endmodule
